interface HA_if;
  logic [3:0]a;
  logic [3:0]b;
  logic [3:0]sum;
  logic carry;
endinterface
